MACRO RIGHT
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN RIGHT 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal1 ;
        RECT 0.00000000 30500.00000000 48000.00000000 33500.00000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal1 ;
        RECT 0.00000000 -1500.00000000 48000.00000000 1500.00000000 ;
    END
  END GND

  PIN OUT_T
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 43000.00000000 8500.00000000 45000.00000000 10500.00000000 ;
    END
  END OUT_T

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 7000.00000000 9500.00000000 9000.00000000 11500.00000000 ;
    END
  END A

  PIN EN
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 23000.00000000 20500.00000000 33000.00000000 22500.00000000 ;
    END
  END EN


END RIGHT
