MACRO MIDDLE
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN MIDDLE 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal1 ;
        RECT 0.00000000 30500.00000000 48000.00000000 33500.00000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal1 ;
        RECT 0.00000000 -1500.00000000 48000.00000000 1500.00000000 ;
    END
  END GND

  PIN PO
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 19000.00000000 8500.00000000 21000.00000000 22500.00000000 ;
    END
  END PO

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 23000.00000000 12500.00000000 25000.00000000 22500.00000000 ;
    END
  END Y

  PIN OUT_T
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 7000.00000000 9500.00000000 9000.00000000 22500.00000000 ;
    END
  END OUT_T

  PIN PI
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 15000.00000000 12500.00000000 17000.00000000 22500.00000000 ;
    END
  END PI


END MIDDLE
