MACRO GPIORIGHT
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN GPIORIGHT 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal1 ;
        RECT 0.00000000 30500.00000000 56000.00000000 33500.00000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal1 ;
        RECT 0.00000000 -1500.00000000 56000.00000000 1500.00000000 ;
    END
  END GND

  PIN OUT_T
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 3000.00000000 8500.00000000 5000.00000000 10500.00000000 ;
    END
  END OUT_T

  PIN EN
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 15000.00000000 8500.00000000 17000.00000000 22500.00000000 ;
    END
  END EN

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 31000.00000000 20500.00000000 33000.00000000 22500.00000000 ;
    END
  END A


END GPIORIGHT
